// LAB4 constants.
`ifndef _LAB4_VH_
 `define _LAB4_VH_

 `define LAB4_WR_WIDTH 5
 `define LAB4_REG_WIDTH 24

`endif
