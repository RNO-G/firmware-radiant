`ifndef RADIANT_DEBUG_VH
 `define RADIANT_DEBUG_VH

 `define LAB4D_SHIFT_REGISTER_DEBUG "FALSE"
 `define RAD_ID_CTRL_SPI_DEBUG "FALSE"
 `define RAD_ID_CTRL_JTAG_DEBUG "TRUE"
 `define WBC_INTERCON_DEBUG "FALSE"
 `define BOARDMAN_INTERFACE_DEBUG "TRUE"
 `define PHASE_SCANNER_DEBUG "TRUE"
 `define RADIANT_TRIG_TOP_DEBUG "TRUE"
`endif
